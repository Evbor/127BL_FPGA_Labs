count_driver_inst : count_driver PORT MAP (
		cin	 => cin_sig,
		clock	 => clock_sig,
		sclr	 => sclr_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);
