const_0_inst : const_0 PORT MAP (
		result	 => result_sig
	);
