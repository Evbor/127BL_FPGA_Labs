BC7_Count_inst : BC7_Count PORT MAP (
		cin	 => cin_sig,
		clock	 => clock_sig,
		sclr	 => sclr_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);
