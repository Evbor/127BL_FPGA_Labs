mf_count1_inst : mf_count1 PORT MAP (
		cin	 => cin_sig,
		clock	 => clock_sig,
		sclr	 => sclr_sig,
		q	 => q_sig
	);
