oscillator_inst : oscillator PORT MAP (
		cin	 => cin_sig,
		clock	 => clock_sig,
		sclr	 => sclr_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);
