mf_const_inst : mf_const PORT MAP (
		result	 => result_sig
	);
