const_4_inst : const_4 PORT MAP (
		result	 => result_sig
	);
