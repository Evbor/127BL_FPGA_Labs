BCD_Count_inst : BCD_Count PORT MAP (
		cin	 => cin_sig,
		clock	 => clock_sig,
		sclr	 => sclr_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);
