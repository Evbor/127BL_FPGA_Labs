// megafunction wizard: %LPM_DECODE%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: LPM_DECODE 

// ============================================================
// File Name: decode.v
// Megafunction Name(s):
// 			LPM_DECODE
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 17.0.0 Build 595 04/25/2017 SJ Standard Edition
// ************************************************************

//Copyright (C) 2017  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel MegaCore Function License Agreement, or other 
//applicable license agreement, including, without limitation, 
//that your use is for the sole purpose of programming logic 
//devices manufactured by Intel and sold by Intel or its 
//authorized distributors.  Please refer to the applicable 
//agreement for further details.

module decode (
	data,
	eq1,
	eq255);

	input	[7:0]  data;
	output	  eq1;
	output	  eq255;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: BaseDec NUMERIC "1"
// Retrieval info: PRIVATE: EnableInput NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: PRIVATE: LPM_PIPELINE NUMERIC "0"
// Retrieval info: PRIVATE: Latency NUMERIC "0"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: aclr NUMERIC "0"
// Retrieval info: PRIVATE: clken NUMERIC "0"
// Retrieval info: PRIVATE: eq0 NUMERIC "0"
// Retrieval info: PRIVATE: eq1 NUMERIC "1"
// Retrieval info: PRIVATE: eq10 NUMERIC "0"
// Retrieval info: PRIVATE: eq100 NUMERIC "0"
// Retrieval info: PRIVATE: eq101 NUMERIC "0"
// Retrieval info: PRIVATE: eq102 NUMERIC "0"
// Retrieval info: PRIVATE: eq103 NUMERIC "0"
// Retrieval info: PRIVATE: eq104 NUMERIC "0"
// Retrieval info: PRIVATE: eq105 NUMERIC "0"
// Retrieval info: PRIVATE: eq106 NUMERIC "0"
// Retrieval info: PRIVATE: eq107 NUMERIC "0"
// Retrieval info: PRIVATE: eq108 NUMERIC "0"
// Retrieval info: PRIVATE: eq109 NUMERIC "0"
// Retrieval info: PRIVATE: eq11 NUMERIC "0"
// Retrieval info: PRIVATE: eq110 NUMERIC "0"
// Retrieval info: PRIVATE: eq111 NUMERIC "0"
// Retrieval info: PRIVATE: eq112 NUMERIC "0"
// Retrieval info: PRIVATE: eq113 NUMERIC "0"
// Retrieval info: PRIVATE: eq114 NUMERIC "0"
// Retrieval info: PRIVATE: eq115 NUMERIC "0"
// Retrieval info: PRIVATE: eq116 NUMERIC "0"
// Retrieval info: PRIVATE: eq117 NUMERIC "0"
// Retrieval info: PRIVATE: eq118 NUMERIC "0"
// Retrieval info: PRIVATE: eq119 NUMERIC "0"
// Retrieval info: PRIVATE: eq12 NUMERIC "0"
// Retrieval info: PRIVATE: eq120 NUMERIC "0"
// Retrieval info: PRIVATE: eq121 NUMERIC "0"
// Retrieval info: PRIVATE: eq122 NUMERIC "0"
// Retrieval info: PRIVATE: eq123 NUMERIC "0"
// Retrieval info: PRIVATE: eq124 NUMERIC "0"
// Retrieval info: PRIVATE: eq125 NUMERIC "0"
// Retrieval info: PRIVATE: eq126 NUMERIC "0"
// Retrieval info: PRIVATE: eq127 NUMERIC "0"
// Retrieval info: PRIVATE: eq128 NUMERIC "0"
// Retrieval info: PRIVATE: eq129 NUMERIC "0"
// Retrieval info: PRIVATE: eq13 NUMERIC "0"
// Retrieval info: PRIVATE: eq130 NUMERIC "0"
// Retrieval info: PRIVATE: eq131 NUMERIC "0"
// Retrieval info: PRIVATE: eq132 NUMERIC "0"
// Retrieval info: PRIVATE: eq133 NUMERIC "0"
// Retrieval info: PRIVATE: eq134 NUMERIC "0"
// Retrieval info: PRIVATE: eq135 NUMERIC "0"
// Retrieval info: PRIVATE: eq136 NUMERIC "0"
// Retrieval info: PRIVATE: eq137 NUMERIC "0"
// Retrieval info: PRIVATE: eq138 NUMERIC "0"
// Retrieval info: PRIVATE: eq139 NUMERIC "0"
// Retrieval info: PRIVATE: eq14 NUMERIC "0"
// Retrieval info: PRIVATE: eq140 NUMERIC "0"
// Retrieval info: PRIVATE: eq141 NUMERIC "0"
// Retrieval info: PRIVATE: eq142 NUMERIC "0"
// Retrieval info: PRIVATE: eq143 NUMERIC "0"
// Retrieval info: PRIVATE: eq144 NUMERIC "0"
// Retrieval info: PRIVATE: eq145 NUMERIC "0"
// Retrieval info: PRIVATE: eq146 NUMERIC "0"
// Retrieval info: PRIVATE: eq147 NUMERIC "0"
// Retrieval info: PRIVATE: eq148 NUMERIC "0"
// Retrieval info: PRIVATE: eq149 NUMERIC "0"
// Retrieval info: PRIVATE: eq15 NUMERIC "0"
// Retrieval info: PRIVATE: eq150 NUMERIC "0"
// Retrieval info: PRIVATE: eq151 NUMERIC "0"
// Retrieval info: PRIVATE: eq152 NUMERIC "0"
// Retrieval info: PRIVATE: eq153 NUMERIC "0"
// Retrieval info: PRIVATE: eq154 NUMERIC "0"
// Retrieval info: PRIVATE: eq155 NUMERIC "0"
// Retrieval info: PRIVATE: eq156 NUMERIC "0"
// Retrieval info: PRIVATE: eq157 NUMERIC "0"
// Retrieval info: PRIVATE: eq158 NUMERIC "0"
// Retrieval info: PRIVATE: eq159 NUMERIC "0"
// Retrieval info: PRIVATE: eq16 NUMERIC "0"
// Retrieval info: PRIVATE: eq160 NUMERIC "0"
// Retrieval info: PRIVATE: eq161 NUMERIC "0"
// Retrieval info: PRIVATE: eq162 NUMERIC "0"
// Retrieval info: PRIVATE: eq163 NUMERIC "0"
// Retrieval info: PRIVATE: eq164 NUMERIC "0"
// Retrieval info: PRIVATE: eq165 NUMERIC "0"
// Retrieval info: PRIVATE: eq166 NUMERIC "0"
// Retrieval info: PRIVATE: eq167 NUMERIC "0"
// Retrieval info: PRIVATE: eq168 NUMERIC "0"
// Retrieval info: PRIVATE: eq169 NUMERIC "0"
// Retrieval info: PRIVATE: eq17 NUMERIC "0"
// Retrieval info: PRIVATE: eq170 NUMERIC "0"
// Retrieval info: PRIVATE: eq171 NUMERIC "0"
// Retrieval info: PRIVATE: eq172 NUMERIC "0"
// Retrieval info: PRIVATE: eq173 NUMERIC "0"
// Retrieval info: PRIVATE: eq174 NUMERIC "0"
// Retrieval info: PRIVATE: eq175 NUMERIC "0"
// Retrieval info: PRIVATE: eq176 NUMERIC "0"
// Retrieval info: PRIVATE: eq177 NUMERIC "0"
// Retrieval info: PRIVATE: eq178 NUMERIC "0"
// Retrieval info: PRIVATE: eq179 NUMERIC "0"
// Retrieval info: PRIVATE: eq18 NUMERIC "0"
// Retrieval info: PRIVATE: eq180 NUMERIC "0"
// Retrieval info: PRIVATE: eq181 NUMERIC "0"
// Retrieval info: PRIVATE: eq182 NUMERIC "0"
// Retrieval info: PRIVATE: eq183 NUMERIC "0"
// Retrieval info: PRIVATE: eq184 NUMERIC "0"
// Retrieval info: PRIVATE: eq185 NUMERIC "0"
// Retrieval info: PRIVATE: eq186 NUMERIC "0"
// Retrieval info: PRIVATE: eq187 NUMERIC "0"
// Retrieval info: PRIVATE: eq188 NUMERIC "0"
// Retrieval info: PRIVATE: eq189 NUMERIC "0"
// Retrieval info: PRIVATE: eq19 NUMERIC "0"
// Retrieval info: PRIVATE: eq190 NUMERIC "0"
// Retrieval info: PRIVATE: eq191 NUMERIC "0"
// Retrieval info: PRIVATE: eq192 NUMERIC "0"
// Retrieval info: PRIVATE: eq193 NUMERIC "0"
// Retrieval info: PRIVATE: eq194 NUMERIC "0"
// Retrieval info: PRIVATE: eq195 NUMERIC "0"
// Retrieval info: PRIVATE: eq196 NUMERIC "0"
// Retrieval info: PRIVATE: eq197 NUMERIC "0"
// Retrieval info: PRIVATE: eq198 NUMERIC "0"
// Retrieval info: PRIVATE: eq199 NUMERIC "0"
// Retrieval info: PRIVATE: eq2 NUMERIC "0"
// Retrieval info: PRIVATE: eq20 NUMERIC "0"
// Retrieval info: PRIVATE: eq200 NUMERIC "0"
// Retrieval info: PRIVATE: eq201 NUMERIC "0"
// Retrieval info: PRIVATE: eq202 NUMERIC "0"
// Retrieval info: PRIVATE: eq203 NUMERIC "0"
// Retrieval info: PRIVATE: eq204 NUMERIC "0"
// Retrieval info: PRIVATE: eq205 NUMERIC "0"
// Retrieval info: PRIVATE: eq206 NUMERIC "0"
// Retrieval info: PRIVATE: eq207 NUMERIC "0"
// Retrieval info: PRIVATE: eq208 NUMERIC "0"
// Retrieval info: PRIVATE: eq209 NUMERIC "0"
// Retrieval info: PRIVATE: eq21 NUMERIC "0"
// Retrieval info: PRIVATE: eq210 NUMERIC "0"
// Retrieval info: PRIVATE: eq211 NUMERIC "0"
// Retrieval info: PRIVATE: eq212 NUMERIC "0"
// Retrieval info: PRIVATE: eq213 NUMERIC "0"
// Retrieval info: PRIVATE: eq214 NUMERIC "0"
// Retrieval info: PRIVATE: eq215 NUMERIC "0"
// Retrieval info: PRIVATE: eq216 NUMERIC "0"
// Retrieval info: PRIVATE: eq217 NUMERIC "0"
// Retrieval info: PRIVATE: eq218 NUMERIC "0"
// Retrieval info: PRIVATE: eq219 NUMERIC "0"
// Retrieval info: PRIVATE: eq22 NUMERIC "0"
// Retrieval info: PRIVATE: eq220 NUMERIC "0"
// Retrieval info: PRIVATE: eq221 NUMERIC "0"
// Retrieval info: PRIVATE: eq222 NUMERIC "0"
// Retrieval info: PRIVATE: eq223 NUMERIC "0"
// Retrieval info: PRIVATE: eq224 NUMERIC "0"
// Retrieval info: PRIVATE: eq225 NUMERIC "0"
// Retrieval info: PRIVATE: eq226 NUMERIC "0"
// Retrieval info: PRIVATE: eq227 NUMERIC "0"
// Retrieval info: PRIVATE: eq228 NUMERIC "0"
// Retrieval info: PRIVATE: eq229 NUMERIC "0"
// Retrieval info: PRIVATE: eq23 NUMERIC "0"
// Retrieval info: PRIVATE: eq230 NUMERIC "0"
// Retrieval info: PRIVATE: eq231 NUMERIC "0"
// Retrieval info: PRIVATE: eq232 NUMERIC "0"
// Retrieval info: PRIVATE: eq233 NUMERIC "0"
// Retrieval info: PRIVATE: eq234 NUMERIC "0"
// Retrieval info: PRIVATE: eq235 NUMERIC "0"
// Retrieval info: PRIVATE: eq236 NUMERIC "0"
// Retrieval info: PRIVATE: eq237 NUMERIC "0"
// Retrieval info: PRIVATE: eq238 NUMERIC "0"
// Retrieval info: PRIVATE: eq239 NUMERIC "0"
// Retrieval info: PRIVATE: eq24 NUMERIC "0"
// Retrieval info: PRIVATE: eq240 NUMERIC "0"
// Retrieval info: PRIVATE: eq241 NUMERIC "0"
// Retrieval info: PRIVATE: eq242 NUMERIC "0"
// Retrieval info: PRIVATE: eq243 NUMERIC "0"
// Retrieval info: PRIVATE: eq244 NUMERIC "0"
// Retrieval info: PRIVATE: eq245 NUMERIC "0"
// Retrieval info: PRIVATE: eq246 NUMERIC "0"
// Retrieval info: PRIVATE: eq247 NUMERIC "0"
// Retrieval info: PRIVATE: eq248 NUMERIC "0"
// Retrieval info: PRIVATE: eq249 NUMERIC "0"
// Retrieval info: PRIVATE: eq25 NUMERIC "0"
// Retrieval info: PRIVATE: eq250 NUMERIC "0"
// Retrieval info: PRIVATE: eq251 NUMERIC "0"
// Retrieval info: PRIVATE: eq252 NUMERIC "0"
// Retrieval info: PRIVATE: eq253 NUMERIC "0"
// Retrieval info: PRIVATE: eq254 NUMERIC "0"
// Retrieval info: PRIVATE: eq255 NUMERIC "1"
// Retrieval info: PRIVATE: eq26 NUMERIC "0"
// Retrieval info: PRIVATE: eq27 NUMERIC "0"
// Retrieval info: PRIVATE: eq28 NUMERIC "0"
// Retrieval info: PRIVATE: eq29 NUMERIC "0"
// Retrieval info: PRIVATE: eq3 NUMERIC "0"
// Retrieval info: PRIVATE: eq30 NUMERIC "0"
// Retrieval info: PRIVATE: eq31 NUMERIC "0"
// Retrieval info: PRIVATE: eq32 NUMERIC "0"
// Retrieval info: PRIVATE: eq33 NUMERIC "0"
// Retrieval info: PRIVATE: eq34 NUMERIC "0"
// Retrieval info: PRIVATE: eq35 NUMERIC "0"
// Retrieval info: PRIVATE: eq36 NUMERIC "0"
// Retrieval info: PRIVATE: eq37 NUMERIC "0"
// Retrieval info: PRIVATE: eq38 NUMERIC "0"
// Retrieval info: PRIVATE: eq39 NUMERIC "0"
// Retrieval info: PRIVATE: eq4 NUMERIC "0"
// Retrieval info: PRIVATE: eq40 NUMERIC "0"
// Retrieval info: PRIVATE: eq41 NUMERIC "0"
// Retrieval info: PRIVATE: eq42 NUMERIC "0"
// Retrieval info: PRIVATE: eq43 NUMERIC "0"
// Retrieval info: PRIVATE: eq44 NUMERIC "0"
// Retrieval info: PRIVATE: eq45 NUMERIC "0"
// Retrieval info: PRIVATE: eq46 NUMERIC "0"
// Retrieval info: PRIVATE: eq47 NUMERIC "0"
// Retrieval info: PRIVATE: eq48 NUMERIC "0"
// Retrieval info: PRIVATE: eq49 NUMERIC "0"
// Retrieval info: PRIVATE: eq5 NUMERIC "0"
// Retrieval info: PRIVATE: eq50 NUMERIC "0"
// Retrieval info: PRIVATE: eq51 NUMERIC "0"
// Retrieval info: PRIVATE: eq52 NUMERIC "0"
// Retrieval info: PRIVATE: eq53 NUMERIC "0"
// Retrieval info: PRIVATE: eq54 NUMERIC "0"
// Retrieval info: PRIVATE: eq55 NUMERIC "0"
// Retrieval info: PRIVATE: eq56 NUMERIC "0"
// Retrieval info: PRIVATE: eq57 NUMERIC "0"
// Retrieval info: PRIVATE: eq58 NUMERIC "0"
// Retrieval info: PRIVATE: eq59 NUMERIC "0"
// Retrieval info: PRIVATE: eq6 NUMERIC "0"
// Retrieval info: PRIVATE: eq60 NUMERIC "0"
// Retrieval info: PRIVATE: eq61 NUMERIC "0"
// Retrieval info: PRIVATE: eq62 NUMERIC "0"
// Retrieval info: PRIVATE: eq63 NUMERIC "0"
// Retrieval info: PRIVATE: eq64 NUMERIC "0"
// Retrieval info: PRIVATE: eq65 NUMERIC "0"
// Retrieval info: PRIVATE: eq66 NUMERIC "0"
// Retrieval info: PRIVATE: eq67 NUMERIC "0"
// Retrieval info: PRIVATE: eq68 NUMERIC "0"
// Retrieval info: PRIVATE: eq69 NUMERIC "0"
// Retrieval info: PRIVATE: eq7 NUMERIC "0"
// Retrieval info: PRIVATE: eq70 NUMERIC "0"
// Retrieval info: PRIVATE: eq71 NUMERIC "0"
// Retrieval info: PRIVATE: eq72 NUMERIC "0"
// Retrieval info: PRIVATE: eq73 NUMERIC "0"
// Retrieval info: PRIVATE: eq74 NUMERIC "0"
// Retrieval info: PRIVATE: eq75 NUMERIC "0"
// Retrieval info: PRIVATE: eq76 NUMERIC "0"
// Retrieval info: PRIVATE: eq77 NUMERIC "0"
// Retrieval info: PRIVATE: eq78 NUMERIC "0"
// Retrieval info: PRIVATE: eq79 NUMERIC "0"
// Retrieval info: PRIVATE: eq8 NUMERIC "0"
// Retrieval info: PRIVATE: eq80 NUMERIC "0"
// Retrieval info: PRIVATE: eq81 NUMERIC "0"
// Retrieval info: PRIVATE: eq82 NUMERIC "0"
// Retrieval info: PRIVATE: eq83 NUMERIC "0"
// Retrieval info: PRIVATE: eq84 NUMERIC "0"
// Retrieval info: PRIVATE: eq85 NUMERIC "0"
// Retrieval info: PRIVATE: eq86 NUMERIC "0"
// Retrieval info: PRIVATE: eq87 NUMERIC "0"
// Retrieval info: PRIVATE: eq88 NUMERIC "0"
// Retrieval info: PRIVATE: eq89 NUMERIC "0"
// Retrieval info: PRIVATE: eq9 NUMERIC "0"
// Retrieval info: PRIVATE: eq90 NUMERIC "0"
// Retrieval info: PRIVATE: eq91 NUMERIC "0"
// Retrieval info: PRIVATE: eq92 NUMERIC "0"
// Retrieval info: PRIVATE: eq93 NUMERIC "0"
// Retrieval info: PRIVATE: eq94 NUMERIC "0"
// Retrieval info: PRIVATE: eq95 NUMERIC "0"
// Retrieval info: PRIVATE: eq96 NUMERIC "0"
// Retrieval info: PRIVATE: eq97 NUMERIC "0"
// Retrieval info: PRIVATE: eq98 NUMERIC "0"
// Retrieval info: PRIVATE: eq99 NUMERIC "0"
// Retrieval info: PRIVATE: nBit NUMERIC "8"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_DECODES NUMERIC "256"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_DECODE"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "8"
// Retrieval info: USED_PORT: @eq 0 0 256 0 OUTPUT NODEFVAL "@eq[255..0]"
// Retrieval info: USED_PORT: data 0 0 8 0 INPUT NODEFVAL "data[7..0]"
// Retrieval info: USED_PORT: eq1 0 0 0 0 OUTPUT NODEFVAL "eq1"
// Retrieval info: USED_PORT: eq255 0 0 0 0 OUTPUT NODEFVAL "eq255"
// Retrieval info: CONNECT: @data 0 0 8 0 data 0 0 8 0
// Retrieval info: CONNECT: eq1 0 0 0 0 @eq 0 0 1 1
// Retrieval info: CONNECT: eq255 0 0 0 0 @eq 0 0 1 255
// Retrieval info: GEN_FILE: TYPE_NORMAL decode.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL decode.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL decode.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL decode.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL decode_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL decode_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
